module MixColumns()