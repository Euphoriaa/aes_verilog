module SubBytes #(parameter numbytes = 16) (input [(8*numbytes - 1):0] in, output reg [(8*numbytes-1):0] out);
    integer i;
    reg [7:0] address;
    always@(*) begin
        for(i = 0; i < numbytes; i = i + 1) begin
            address = in[i*8 +: 8];
            case (address)
                8'h0 : out[i*8+:8] = 8'h63;
                8'h1 : out[i*8+:8] = 8'h7C;
                8'h2 : out[i*8+:8] = 8'h77;
                8'h3 : out[i*8+:8] = 8'h7B;
                8'h4 : out[i*8+:8] = 8'hF2;
                8'h5 : out[i*8+:8] = 8'h6B;
                8'h6 : out[i*8+:8] = 8'h6F;
                8'h7 : out[i*8+:8] = 8'hC5;
                8'h8 : out[i*8+:8] = 8'h30;
                8'h9 : out[i*8+:8] = 8'h1;
                8'hA : out[i*8+:8] = 8'h67;
                8'hB : out[i*8+:8] = 8'h2B;
                8'hC : out[i*8+:8] = 8'hFE;
                8'hD : out[i*8+:8] = 8'hD7;
                8'hE : out[i*8+:8] = 8'hAB;
                8'hF : out[i*8+:8] = 8'h76;
                8'h10 : out[i*8+:8] = 8'hCA;
                8'h11 : out[i*8+:8] = 8'h82;
                8'h12 : out[i*8+:8] = 8'hC9;
                8'h13 : out[i*8+:8] = 8'h7D;
                8'h14 : out[i*8+:8] = 8'hFA;
                8'h15 : out[i*8+:8] = 8'h59;
                8'h16 : out[i*8+:8] = 8'h47;
                8'h17 : out[i*8+:8] = 8'hF0;
                8'h18 : out[i*8+:8] = 8'hAD;
                8'h19 : out[i*8+:8] = 8'hD4;
                8'h1A : out[i*8+:8] = 8'hA2;
                8'h1B : out[i*8+:8] = 8'hAF;
                8'h1C : out[i*8+:8] = 8'h9C;
                8'h1D : out[i*8+:8] = 8'hA4;
                8'h1E : out[i*8+:8] = 8'h72;
                8'h1F : out[i*8+:8] = 8'hC0;
                8'h20 : out[i*8+:8] = 8'hB7;
                8'h21 : out[i*8+:8] = 8'hFD;
                8'h22 : out[i*8+:8] = 8'h93;
                8'h23 : out[i*8+:8] = 8'h26;
                8'h24 : out[i*8+:8] = 8'h36;
                8'h25 : out[i*8+:8] = 8'h3F;
                8'h26 : out[i*8+:8] = 8'hF7;
                8'h27 : out[i*8+:8] = 8'hCC;
                8'h28 : out[i*8+:8] = 8'h34;
                8'h29 : out[i*8+:8] = 8'hA5;
                8'h2A : out[i*8+:8] = 8'hE5;
                8'h2B : out[i*8+:8] = 8'hF1;
                8'h2C : out[i*8+:8] = 8'h71;
                8'h2D : out[i*8+:8] = 8'hD8;
                8'h2E : out[i*8+:8] = 8'h31;
                8'h2F : out[i*8+:8] = 8'h15;
                8'h30 : out[i*8+:8] = 8'h4;
                8'h31 : out[i*8+:8] = 8'hC7;
                8'h32 : out[i*8+:8] = 8'h23;
                8'h33 : out[i*8+:8] = 8'hC3;
                8'h34 : out[i*8+:8] = 8'h18;
                8'h35 : out[i*8+:8] = 8'h96;
                8'h36 : out[i*8+:8] = 8'h5;
                8'h37 : out[i*8+:8] = 8'h9A;
                8'h38 : out[i*8+:8] = 8'h7;
                8'h39 : out[i*8+:8] = 8'h12;
                8'h3A : out[i*8+:8] = 8'h80;
                8'h3B : out[i*8+:8] = 8'hE2;
                8'h3C : out[i*8+:8] = 8'hEB;
                8'h3D : out[i*8+:8] = 8'h27;
                8'h3E : out[i*8+:8] = 8'hB2;
                8'h3F : out[i*8+:8] = 8'h75;
                8'h40 : out[i*8+:8] = 8'h9;
                8'h41 : out[i*8+:8] = 8'h83;
                8'h42 : out[i*8+:8] = 8'h2C;
                8'h43 : out[i*8+:8] = 8'h1A;
                8'h44 : out[i*8+:8] = 8'h1B;
                8'h45 : out[i*8+:8] = 8'h6E;
                8'h46 : out[i*8+:8] = 8'h5A;
                8'h47 : out[i*8+:8] = 8'hA0;
                8'h48 : out[i*8+:8] = 8'h52;
                8'h49 : out[i*8+:8] = 8'h3B;
                8'h4A : out[i*8+:8] = 8'hD6;
                8'h4B : out[i*8+:8] = 8'hB3;
                8'h4C : out[i*8+:8] = 8'h29;
                8'h4D : out[i*8+:8] = 8'hE3;
                8'h4E : out[i*8+:8] = 8'h2F;
                8'h4F : out[i*8+:8] = 8'h84;
                8'h50 : out[i*8+:8] = 8'h53;
                8'h51 : out[i*8+:8] = 8'hD1;
                8'h52 : out[i*8+:8] = 8'h0;
                8'h53 : out[i*8+:8] = 8'hED;
                8'h54 : out[i*8+:8] = 8'h20;
                8'h55 : out[i*8+:8] = 8'hFC;
                8'h56 : out[i*8+:8] = 8'hB1;
                8'h57 : out[i*8+:8] = 8'h5B;
                8'h58 : out[i*8+:8] = 8'h6A;
                8'h59 : out[i*8+:8] = 8'hCB;
                8'h5A : out[i*8+:8] = 8'hBE;
                8'h5B : out[i*8+:8] = 8'h39;
                8'h5C : out[i*8+:8] = 8'h4A;
                8'h5D : out[i*8+:8] = 8'h4C;
                8'h5E : out[i*8+:8] = 8'h58;
                8'h5F : out[i*8+:8] = 8'hCF;
                8'h60 : out[i*8+:8] = 8'hD0;
                8'h61 : out[i*8+:8] = 8'hEF;
                8'h62 : out[i*8+:8] = 8'hAA;
                8'h63 : out[i*8+:8] = 8'hFB;
                8'h64 : out[i*8+:8] = 8'h43;
                8'h65 : out[i*8+:8] = 8'h4D;
                8'h66 : out[i*8+:8] = 8'h33;
                8'h67 : out[i*8+:8] = 8'h85;
                8'h68 : out[i*8+:8] = 8'h45;
                8'h69 : out[i*8+:8] = 8'hF9;
                8'h6A : out[i*8+:8] = 8'h2;
                8'h6B : out[i*8+:8] = 8'h7F;
                8'h6C : out[i*8+:8] = 8'h50;
                8'h6D : out[i*8+:8] = 8'h3C;
                8'h6E : out[i*8+:8] = 8'h9F;
                8'h6F : out[i*8+:8] = 8'hA8;
                8'h70 : out[i*8+:8] = 8'h51;
                8'h71 : out[i*8+:8] = 8'hA3;
                8'h72 : out[i*8+:8] = 8'h40;
                8'h73 : out[i*8+:8] = 8'h8F;
                8'h74 : out[i*8+:8] = 8'h92;
                8'h75 : out[i*8+:8] = 8'h9D;
                8'h76 : out[i*8+:8] = 8'h38;
                8'h77 : out[i*8+:8] = 8'hF5;
                8'h78 : out[i*8+:8] = 8'hBC;
                8'h79 : out[i*8+:8] = 8'hB6;
                8'h7A : out[i*8+:8] = 8'hDA;
                8'h7B : out[i*8+:8] = 8'h21;
                8'h7C : out[i*8+:8] = 8'h10;
                8'h7D : out[i*8+:8] = 8'hFF;
                8'h7E : out[i*8+:8] = 8'hF3;
                8'h7F : out[i*8+:8] = 8'hD2;
                8'h80 : out[i*8+:8] = 8'hCD;
                8'h81 : out[i*8+:8] = 8'hC;
                8'h82 : out[i*8+:8] = 8'h13;
                8'h83 : out[i*8+:8] = 8'hEC;
                8'h84 : out[i*8+:8] = 8'h5F;
                8'h85 : out[i*8+:8] = 8'h97;
                8'h86 : out[i*8+:8] = 8'h44;
                8'h87 : out[i*8+:8] = 8'h17;
                8'h88 : out[i*8+:8] = 8'hC4;
                8'h89 : out[i*8+:8] = 8'hA7;
                8'h8A : out[i*8+:8] = 8'h7E;
                8'h8B : out[i*8+:8] = 8'h3D;
                8'h8C : out[i*8+:8] = 8'h64;
                8'h8D : out[i*8+:8] = 8'h5D;
                8'h8E : out[i*8+:8] = 8'h19;
                8'h8F : out[i*8+:8] = 8'h73;
                8'h90 : out[i*8+:8] = 8'h60;
                8'h91 : out[i*8+:8] = 8'h81;
                8'h92 : out[i*8+:8] = 8'h4F;
                8'h93 : out[i*8+:8] = 8'hDC;
                8'h94 : out[i*8+:8] = 8'h22;
                8'h95 : out[i*8+:8] = 8'h2A;
                8'h96 : out[i*8+:8] = 8'h90;
                8'h97 : out[i*8+:8] = 8'h88;
                8'h98 : out[i*8+:8] = 8'h46;
                8'h99 : out[i*8+:8] = 8'hEE;
                8'h9A : out[i*8+:8] = 8'hB8;
                8'h9B : out[i*8+:8] = 8'h14;
                8'h9C : out[i*8+:8] = 8'hDE;
                8'h9D : out[i*8+:8] = 8'h5E;
                8'h9E : out[i*8+:8] = 8'hB;
                8'h9F : out[i*8+:8] = 8'hDB;
                8'hA0 : out[i*8+:8] = 8'hE0;
                8'hA1 : out[i*8+:8] = 8'h32;
                8'hA2 : out[i*8+:8] = 8'h3A;
                8'hA3 : out[i*8+:8] = 8'hA;
                8'hA4 : out[i*8+:8] = 8'h49;
                8'hA5 : out[i*8+:8] = 8'h6;
                8'hA6 : out[i*8+:8] = 8'h24;
                8'hA7 : out[i*8+:8] = 8'h5C;
                8'hA8 : out[i*8+:8] = 8'hC2;
                8'hA9 : out[i*8+:8] = 8'hD3;
                8'hAA : out[i*8+:8] = 8'hAC;
                8'hAB : out[i*8+:8] = 8'h62;
                8'hAC : out[i*8+:8] = 8'h91;
                8'hAD : out[i*8+:8] = 8'h95;
                8'hAE : out[i*8+:8] = 8'hE4;
                8'hAF : out[i*8+:8] = 8'h79;
                8'hB0 : out[i*8+:8] = 8'hE7;
                8'hB1 : out[i*8+:8] = 8'hC8;
                8'hB2 : out[i*8+:8] = 8'h37;
                8'hB3 : out[i*8+:8] = 8'h6D;
                8'hB4 : out[i*8+:8] = 8'h8D;
                8'hB5 : out[i*8+:8] = 8'hD5;
                8'hB6 : out[i*8+:8] = 8'h4E;
                8'hB7 : out[i*8+:8] = 8'hA9;
                8'hB8 : out[i*8+:8] = 8'h6C;
                8'hB9 : out[i*8+:8] = 8'h56;
                8'hBA : out[i*8+:8] = 8'hF4;
                8'hBB : out[i*8+:8] = 8'hEA;
                8'hBC : out[i*8+:8] = 8'h65;
                8'hBD : out[i*8+:8] = 8'h7A;
                8'hBE : out[i*8+:8] = 8'hAE;
                8'hBF : out[i*8+:8] = 8'h8;
                8'hC0 : out[i*8+:8] = 8'hBA;
                8'hC1 : out[i*8+:8] = 8'h78;
                8'hC2 : out[i*8+:8] = 8'h25;
                8'hC3 : out[i*8+:8] = 8'h2E;
                8'hC4 : out[i*8+:8] = 8'h1C;
                8'hC5 : out[i*8+:8] = 8'hA6;
                8'hC6 : out[i*8+:8] = 8'hB4;
                8'hC7 : out[i*8+:8] = 8'hC6;
                8'hC8 : out[i*8+:8] = 8'hE8;
                8'hC9 : out[i*8+:8] = 8'hDD;
                8'hCA : out[i*8+:8] = 8'h74;
                8'hCB : out[i*8+:8] = 8'h1F;
                8'hCC : out[i*8+:8] = 8'h4B;
                8'hCD : out[i*8+:8] = 8'hBD;
                8'hCE : out[i*8+:8] = 8'h8B;
                8'hCF : out[i*8+:8] = 8'h8A;
                8'hD0 : out[i*8+:8] = 8'h70;
                8'hD1 : out[i*8+:8] = 8'h3E;
                8'hD2 : out[i*8+:8] = 8'hB5;
                8'hD3 : out[i*8+:8] = 8'h66;
                8'hD4 : out[i*8+:8] = 8'h48;
                8'hD5 : out[i*8+:8] = 8'h3;
                8'hD6 : out[i*8+:8] = 8'hF6;
                8'hD7 : out[i*8+:8] = 8'hE;
                8'hD8 : out[i*8+:8] = 8'h61;
                8'hD9 : out[i*8+:8] = 8'h35;
                8'hDA : out[i*8+:8] = 8'h57;
                8'hDB : out[i*8+:8] = 8'hB9;
                8'hDC : out[i*8+:8] = 8'h86;
                8'hDD : out[i*8+:8] = 8'hC1;
                8'hDE : out[i*8+:8] = 8'h1D;
                8'hDF : out[i*8+:8] = 8'h9E;
                8'hE0 : out[i*8+:8] = 8'hE1;
                8'hE1 : out[i*8+:8] = 8'hF8;
                8'hE2 : out[i*8+:8] = 8'h98;
                8'hE3 : out[i*8+:8] = 8'h11;
                8'hE4 : out[i*8+:8] = 8'h69;
                8'hE5 : out[i*8+:8] = 8'hD9;
                8'hE6 : out[i*8+:8] = 8'h8E;
                8'hE7 : out[i*8+:8] = 8'h94;
                8'hE8 : out[i*8+:8] = 8'h9B;
                8'hE9 : out[i*8+:8] = 8'h1E;
                8'hEA : out[i*8+:8] = 8'h87;
                8'hEB : out[i*8+:8] = 8'hE9;
                8'hEC : out[i*8+:8] = 8'hCE;
                8'hED : out[i*8+:8] = 8'h55;
                8'hEE : out[i*8+:8] = 8'h28;
                8'hEF : out[i*8+:8] = 8'hDF;
                8'hF0 : out[i*8+:8] = 8'h8C;
                8'hF1 : out[i*8+:8] = 8'hA1;
                8'hF2 : out[i*8+:8] = 8'h89;
                8'hF3 : out[i*8+:8] = 8'hD;
                8'hF4 : out[i*8+:8] = 8'hBF;
                8'hF5 : out[i*8+:8] = 8'hE6;
                8'hF6 : out[i*8+:8] = 8'h42;
                8'hF7 : out[i*8+:8] = 8'h68;
                8'hF8 : out[i*8+:8] = 8'h41;
                8'hF9 : out[i*8+:8] = 8'h99;
                8'hFA : out[i*8+:8] = 8'h2D;
                8'hFB : out[i*8+:8] = 8'hF;
                8'hFC : out[i*8+:8] = 8'hB0;
                8'hFD : out[i*8+:8] = 8'h54;
                8'hFE : out[i*8+:8] = 8'hBB;
                8'hFF : out[i*8+:8] = 8'h16;
                default : out[i*8+:8] = 8'h0;
            endcase
        end
    end
endmodule