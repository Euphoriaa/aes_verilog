module SubBytes(input [127:0] state, output reg [127:0] nstate);
    integer i;
    reg [7:0] address;
    always@(*) begin
        for(i = 0; i < 16; i = i + 1) begin
            address = state[i*8 +: 8];
            case (address)
                8'h0 : nstate[i*8+:8] = 8'h63;
                8'h1 : nstate[i*8+:8] = 8'h7C;
                8'h2 : nstate[i*8+:8] = 8'h77;
                8'h3 : nstate[i*8+:8] = 8'h7B;
                8'h4 : nstate[i*8+:8] = 8'hF2;
                8'h5 : nstate[i*8+:8] = 8'h6B;
                8'h6 : nstate[i*8+:8] = 8'h6F;
                8'h7 : nstate[i*8+:8] = 8'hC5;
                8'h8 : nstate[i*8+:8] = 8'h30;
                8'h9 : nstate[i*8+:8] = 8'h1;
                8'hA : nstate[i*8+:8] = 8'h67;
                8'hB : nstate[i*8+:8] = 8'h2B;
                8'hC : nstate[i*8+:8] = 8'hFE;
                8'hD : nstate[i*8+:8] = 8'hD7;
                8'hE : nstate[i*8+:8] = 8'hAB;
                8'hF : nstate[i*8+:8] = 8'h76;
                8'h10 : nstate[i*8+:8] = 8'hCA;
                8'h11 : nstate[i*8+:8] = 8'h82;
                8'h12 : nstate[i*8+:8] = 8'hC9;
                8'h13 : nstate[i*8+:8] = 8'h7D;
                8'h14 : nstate[i*8+:8] = 8'hFA;
                8'h15 : nstate[i*8+:8] = 8'h59;
                8'h16 : nstate[i*8+:8] = 8'h47;
                8'h17 : nstate[i*8+:8] = 8'hF0;
                8'h18 : nstate[i*8+:8] = 8'hAD;
                8'h19 : nstate[i*8+:8] = 8'hD4;
                8'h1A : nstate[i*8+:8] = 8'hA2;
                8'h1B : nstate[i*8+:8] = 8'hAF;
                8'h1C : nstate[i*8+:8] = 8'h9C;
                8'h1D : nstate[i*8+:8] = 8'hA4;
                8'h1E : nstate[i*8+:8] = 8'h72;
                8'h1F : nstate[i*8+:8] = 8'hC0;
                8'h20 : nstate[i*8+:8] = 8'hB7;
                8'h21 : nstate[i*8+:8] = 8'hFD;
                8'h22 : nstate[i*8+:8] = 8'h93;
                8'h23 : nstate[i*8+:8] = 8'h26;
                8'h24 : nstate[i*8+:8] = 8'h36;
                8'h25 : nstate[i*8+:8] = 8'h3F;
                8'h26 : nstate[i*8+:8] = 8'hF7;
                8'h27 : nstate[i*8+:8] = 8'hCC;
                8'h28 : nstate[i*8+:8] = 8'h34;
                8'h29 : nstate[i*8+:8] = 8'hA5;
                8'h2A : nstate[i*8+:8] = 8'hE5;
                8'h2B : nstate[i*8+:8] = 8'hF1;
                8'h2C : nstate[i*8+:8] = 8'h71;
                8'h2D : nstate[i*8+:8] = 8'hD8;
                8'h2E : nstate[i*8+:8] = 8'h31;
                8'h2F : nstate[i*8+:8] = 8'h15;
                8'h30 : nstate[i*8+:8] = 8'h4;
                8'h31 : nstate[i*8+:8] = 8'hC7;
                8'h32 : nstate[i*8+:8] = 8'h23;
                8'h33 : nstate[i*8+:8] = 8'hC3;
                8'h34 : nstate[i*8+:8] = 8'h18;
                8'h35 : nstate[i*8+:8] = 8'h96;
                8'h36 : nstate[i*8+:8] = 8'h5;
                8'h37 : nstate[i*8+:8] = 8'h9A;
                8'h38 : nstate[i*8+:8] = 8'h7;
                8'h39 : nstate[i*8+:8] = 8'h12;
                8'h3A : nstate[i*8+:8] = 8'h80;
                8'h3B : nstate[i*8+:8] = 8'hE2;
                8'h3C : nstate[i*8+:8] = 8'hEB;
                8'h3D : nstate[i*8+:8] = 8'h27;
                8'h3E : nstate[i*8+:8] = 8'hB2;
                8'h3F : nstate[i*8+:8] = 8'h75;
                8'h40 : nstate[i*8+:8] = 8'h9;
                8'h41 : nstate[i*8+:8] = 8'h83;
                8'h42 : nstate[i*8+:8] = 8'h2C;
                8'h43 : nstate[i*8+:8] = 8'h1A;
                8'h44 : nstate[i*8+:8] = 8'h1B;
                8'h45 : nstate[i*8+:8] = 8'h6E;
                8'h46 : nstate[i*8+:8] = 8'h5A;
                8'h47 : nstate[i*8+:8] = 8'hA0;
                8'h48 : nstate[i*8+:8] = 8'h52;
                8'h49 : nstate[i*8+:8] = 8'h3B;
                8'h4A : nstate[i*8+:8] = 8'hD6;
                8'h4B : nstate[i*8+:8] = 8'hB3;
                8'h4C : nstate[i*8+:8] = 8'h29;
                8'h4D : nstate[i*8+:8] = 8'hE3;
                8'h4E : nstate[i*8+:8] = 8'h2F;
                8'h4F : nstate[i*8+:8] = 8'h84;
                8'h50 : nstate[i*8+:8] = 8'h53;
                8'h51 : nstate[i*8+:8] = 8'hD1;
                8'h52 : nstate[i*8+:8] = 8'h0;
                8'h53 : nstate[i*8+:8] = 8'hED;
                8'h54 : nstate[i*8+:8] = 8'h20;
                8'h55 : nstate[i*8+:8] = 8'hFC;
                8'h56 : nstate[i*8+:8] = 8'hB1;
                8'h57 : nstate[i*8+:8] = 8'h5B;
                8'h58 : nstate[i*8+:8] = 8'h6A;
                8'h59 : nstate[i*8+:8] = 8'hCB;
                8'h5A : nstate[i*8+:8] = 8'hBE;
                8'h5B : nstate[i*8+:8] = 8'h39;
                8'h5C : nstate[i*8+:8] = 8'h4A;
                8'h5D : nstate[i*8+:8] = 8'h4C;
                8'h5E : nstate[i*8+:8] = 8'h58;
                8'h5F : nstate[i*8+:8] = 8'hCF;
                8'h60 : nstate[i*8+:8] = 8'hD0;
                8'h61 : nstate[i*8+:8] = 8'hEF;
                8'h62 : nstate[i*8+:8] = 8'hAA;
                8'h63 : nstate[i*8+:8] = 8'hFB;
                8'h64 : nstate[i*8+:8] = 8'h43;
                8'h65 : nstate[i*8+:8] = 8'h4D;
                8'h66 : nstate[i*8+:8] = 8'h33;
                8'h67 : nstate[i*8+:8] = 8'h85;
                8'h68 : nstate[i*8+:8] = 8'h45;
                8'h69 : nstate[i*8+:8] = 8'hF9;
                8'h6A : nstate[i*8+:8] = 8'h2;
                8'h6B : nstate[i*8+:8] = 8'h7F;
                8'h6C : nstate[i*8+:8] = 8'h50;
                8'h6D : nstate[i*8+:8] = 8'h3C;
                8'h6E : nstate[i*8+:8] = 8'h9F;
                8'h6F : nstate[i*8+:8] = 8'hA8;
                8'h70 : nstate[i*8+:8] = 8'h51;
                8'h71 : nstate[i*8+:8] = 8'hA3;
                8'h72 : nstate[i*8+:8] = 8'h40;
                8'h73 : nstate[i*8+:8] = 8'h8F;
                8'h74 : nstate[i*8+:8] = 8'h92;
                8'h75 : nstate[i*8+:8] = 8'h9D;
                8'h76 : nstate[i*8+:8] = 8'h38;
                8'h77 : nstate[i*8+:8] = 8'hF5;
                8'h78 : nstate[i*8+:8] = 8'hBC;
                8'h79 : nstate[i*8+:8] = 8'hB6;
                8'h7A : nstate[i*8+:8] = 8'hDA;
                8'h7B : nstate[i*8+:8] = 8'h21;
                8'h7C : nstate[i*8+:8] = 8'h10;
                8'h7D : nstate[i*8+:8] = 8'hFF;
                8'h7E : nstate[i*8+:8] = 8'hF3;
                8'h7F : nstate[i*8+:8] = 8'hD2;
                8'h80 : nstate[i*8+:8] = 8'hCD;
                8'h81 : nstate[i*8+:8] = 8'hC;
                8'h82 : nstate[i*8+:8] = 8'h13;
                8'h83 : nstate[i*8+:8] = 8'hEC;
                8'h84 : nstate[i*8+:8] = 8'h5F;
                8'h85 : nstate[i*8+:8] = 8'h97;
                8'h86 : nstate[i*8+:8] = 8'h44;
                8'h87 : nstate[i*8+:8] = 8'h17;
                8'h88 : nstate[i*8+:8] = 8'hC4;
                8'h89 : nstate[i*8+:8] = 8'hA7;
                8'h8A : nstate[i*8+:8] = 8'h7E;
                8'h8B : nstate[i*8+:8] = 8'h3D;
                8'h8C : nstate[i*8+:8] = 8'h64;
                8'h8D : nstate[i*8+:8] = 8'h5D;
                8'h8E : nstate[i*8+:8] = 8'h19;
                8'h8F : nstate[i*8+:8] = 8'h73;
                8'h90 : nstate[i*8+:8] = 8'h60;
                8'h91 : nstate[i*8+:8] = 8'h81;
                8'h92 : nstate[i*8+:8] = 8'h4F;
                8'h93 : nstate[i*8+:8] = 8'hDC;
                8'h94 : nstate[i*8+:8] = 8'h22;
                8'h95 : nstate[i*8+:8] = 8'h2A;
                8'h96 : nstate[i*8+:8] = 8'h90;
                8'h97 : nstate[i*8+:8] = 8'h88;
                8'h98 : nstate[i*8+:8] = 8'h46;
                8'h99 : nstate[i*8+:8] = 8'hEE;
                8'h9A : nstate[i*8+:8] = 8'hB8;
                8'h9B : nstate[i*8+:8] = 8'h14;
                8'h9C : nstate[i*8+:8] = 8'hDE;
                8'h9D : nstate[i*8+:8] = 8'h5E;
                8'h9E : nstate[i*8+:8] = 8'hB;
                8'h9F : nstate[i*8+:8] = 8'hDB;
                8'hA0 : nstate[i*8+:8] = 8'hE0;
                8'hA1 : nstate[i*8+:8] = 8'h32;
                8'hA2 : nstate[i*8+:8] = 8'h3A;
                8'hA3 : nstate[i*8+:8] = 8'hA;
                8'hA4 : nstate[i*8+:8] = 8'h49;
                8'hA5 : nstate[i*8+:8] = 8'h6;
                8'hA6 : nstate[i*8+:8] = 8'h24;
                8'hA7 : nstate[i*8+:8] = 8'h5C;
                8'hA8 : nstate[i*8+:8] = 8'hC2;
                8'hA9 : nstate[i*8+:8] = 8'hD3;
                8'hAA : nstate[i*8+:8] = 8'hAC;
                8'hAB : nstate[i*8+:8] = 8'h62;
                8'hAC : nstate[i*8+:8] = 8'h91;
                8'hAD : nstate[i*8+:8] = 8'h95;
                8'hAE : nstate[i*8+:8] = 8'hE4;
                8'hAF : nstate[i*8+:8] = 8'h79;
                8'hB0 : nstate[i*8+:8] = 8'hE7;
                8'hB1 : nstate[i*8+:8] = 8'hC8;
                8'hB2 : nstate[i*8+:8] = 8'h37;
                8'hB3 : nstate[i*8+:8] = 8'h6D;
                8'hB4 : nstate[i*8+:8] = 8'h8D;
                8'hB5 : nstate[i*8+:8] = 8'hD5;
                8'hB6 : nstate[i*8+:8] = 8'h4E;
                8'hB7 : nstate[i*8+:8] = 8'hA9;
                8'hB8 : nstate[i*8+:8] = 8'h6C;
                8'hB9 : nstate[i*8+:8] = 8'h56;
                8'hBA : nstate[i*8+:8] = 8'hF4;
                8'hBB : nstate[i*8+:8] = 8'hEA;
                8'hBC : nstate[i*8+:8] = 8'h65;
                8'hBD : nstate[i*8+:8] = 8'h7A;
                8'hBE : nstate[i*8+:8] = 8'hAE;
                8'hBF : nstate[i*8+:8] = 8'h8;
                8'hC0 : nstate[i*8+:8] = 8'hBA;
                8'hC1 : nstate[i*8+:8] = 8'h78;
                8'hC2 : nstate[i*8+:8] = 8'h25;
                8'hC3 : nstate[i*8+:8] = 8'h2E;
                8'hC4 : nstate[i*8+:8] = 8'h1C;
                8'hC5 : nstate[i*8+:8] = 8'hA6;
                8'hC6 : nstate[i*8+:8] = 8'hB4;
                8'hC7 : nstate[i*8+:8] = 8'hC6;
                8'hC8 : nstate[i*8+:8] = 8'hE8;
                8'hC9 : nstate[i*8+:8] = 8'hDD;
                8'hCA : nstate[i*8+:8] = 8'h74;
                8'hCB : nstate[i*8+:8] = 8'h1F;
                8'hCC : nstate[i*8+:8] = 8'h4B;
                8'hCD : nstate[i*8+:8] = 8'hBD;
                8'hCE : nstate[i*8+:8] = 8'h8B;
                8'hCF : nstate[i*8+:8] = 8'h8A;
                8'hD0 : nstate[i*8+:8] = 8'h70;
                8'hD1 : nstate[i*8+:8] = 8'h3E;
                8'hD2 : nstate[i*8+:8] = 8'hB5;
                8'hD3 : nstate[i*8+:8] = 8'h66;
                8'hD4 : nstate[i*8+:8] = 8'h48;
                8'hD5 : nstate[i*8+:8] = 8'h3;
                8'hD6 : nstate[i*8+:8] = 8'hF6;
                8'hD7 : nstate[i*8+:8] = 8'hE;
                8'hD8 : nstate[i*8+:8] = 8'h61;
                8'hD9 : nstate[i*8+:8] = 8'h35;
                8'hDA : nstate[i*8+:8] = 8'h57;
                8'hDB : nstate[i*8+:8] = 8'hB9;
                8'hDC : nstate[i*8+:8] = 8'h86;
                8'hDD : nstate[i*8+:8] = 8'hC1;
                8'hDE : nstate[i*8+:8] = 8'h1D;
                8'hDF : nstate[i*8+:8] = 8'h9E;
                8'hE0 : nstate[i*8+:8] = 8'hE1;
                8'hE1 : nstate[i*8+:8] = 8'hF8;
                8'hE2 : nstate[i*8+:8] = 8'h98;
                8'hE3 : nstate[i*8+:8] = 8'h11;
                8'hE4 : nstate[i*8+:8] = 8'h69;
                8'hE5 : nstate[i*8+:8] = 8'hD9;
                8'hE6 : nstate[i*8+:8] = 8'h8E;
                8'hE7 : nstate[i*8+:8] = 8'h94;
                8'hE8 : nstate[i*8+:8] = 8'h9B;
                8'hE9 : nstate[i*8+:8] = 8'h1E;
                8'hEA : nstate[i*8+:8] = 8'h87;
                8'hEB : nstate[i*8+:8] = 8'hE9;
                8'hEC : nstate[i*8+:8] = 8'hCE;
                8'hED : nstate[i*8+:8] = 8'h55;
                8'hEE : nstate[i*8+:8] = 8'h28;
                8'hEF : nstate[i*8+:8] = 8'hDF;
                8'hF0 : nstate[i*8+:8] = 8'h8C;
                8'hF1 : nstate[i*8+:8] = 8'hA1;
                8'hF2 : nstate[i*8+:8] = 8'h89;
                8'hF3 : nstate[i*8+:8] = 8'hD;
                8'hF4 : nstate[i*8+:8] = 8'hBF;
                8'hF5 : nstate[i*8+:8] = 8'hE6;
                8'hF6 : nstate[i*8+:8] = 8'h42;
                8'hF7 : nstate[i*8+:8] = 8'h68;
                8'hF8 : nstate[i*8+:8] = 8'h41;
                8'hF9 : nstate[i*8+:8] = 8'h99;
                8'hFA : nstate[i*8+:8] = 8'h2D;
                8'hFB : nstate[i*8+:8] = 8'hF;
                8'hFC : nstate[i*8+:8] = 8'hB0;
                8'hFD : nstate[i*8+:8] = 8'h54;
                8'hFE : nstate[i*8+:8] = 8'hBB;
                8'hFF : nstate[i*8+:8] = 8'h16;
                default : nstate[i*8+:8] = 8'h0;
            endcase
        end
    end
endmodule